`timescale 1ns / 1ps

module tb_clock_gated_approx_mult_8bit;

    reg clk;
    reg rst;
    reg en;
    reg [7:0] A, B;
    wire [15:0] Y;

    // DUT
    clock_gated_approx_mult_8bit DUT (
        .clk(clk),
        .rst(rst),
        .en(en),
        .A(A),
        .B(B),
        .Y(Y)
    );

    // Clock generation
    always #5 clk = ~clk;

    initial begin
        clk = 0;
        rst = 1;
        en  = 0;
        A   = 0;
        B   = 0;

        #10 rst = 0;

        // Enable ON → output updates
        en = 1;
        A = 8'd5;   B = 8'd3;    #10;   // ~15
        A = 8'd12;  B = 8'd7;    #10;   // ~84
        A = 8'd25;  B = 8'd4;    #10;   // ~100
        A = 8'd50;  B = 8'd10;   #10;   // ~500

        // Disable → output should HOLD
        en = 0;
        A = 8'd200; B = 8'd200;  #20;
        A = 8'd255; B = 8'd255;  #20;

        // Enable again
        en = 1;
        A = 8'd15;  B = 8'd15;   #10;

        $finish;
    end

endmodule
